library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity and_gate is
   generic (N: integer:= 32);
   port(in1,in2: in std_logic_vector(N-1 downto 0);
        out1      : out std_logic_vector(N-1 downto 0));
end and_gate;

architecture behavioral of and_gate is
   signal  gate1 : std_logic_vector(N-1 downto 0);
begin
   process(in1,in2,gate1)
	   begin
		   for I in 0 to N-1 loop
		     if    in2(I)='0' then gate1(I)<='0';
			  elsif in2(I)='1' then gate1(I)<= in1(I);
			  else  gate1(I)<='X';
			  end if;
		     out1(I)<= gate1(I);
		   end loop;
	end process;
end behavioral;