library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity nand_gate is
   generic (N: integer:= 32);
   port(in1,in2: in std_logic_vector(N-1 downto 0);
        out2      : out std_logic_vector(N-1 downto 0));
end nand_gate;

architecture behavioral of nand_gate is
   signal  gate2 : std_logic_vector(N-1 downto 0);
begin
   process(in1,in2,gate2)
	   begin
		   for I in 0 to N-1 loop
		     if    in2(I)='0' then gate2(I)<=not in2(I);
			  elsif in2(I)='1' then gate2(I)<=not in1(I);
			  else  gate2(I)<='X';
			  end if;
		     out2(I)<= gate2(I);
		   end loop;
	end process;
end behavioral;